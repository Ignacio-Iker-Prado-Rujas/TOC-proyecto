------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : pokemonpeque.ppm 
--- Filas    : 256 
--- Columnas : 256 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_pokemonpeque is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(16-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_pokemonpeque;


architecture BEHAVIORAL of ROM_RGB_9b_pokemonpeque is
  signal addr_int  : natural range 0 to 2**16-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "010010010",
       "001001001",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "001001001",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "000000000",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "000000001",
       "001001010",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000001001",
       "010010010",
       "001001010",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "001001001",
       "000000000",
       "001001001",
       "010010010",
       "001010010",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "001001001",
       "000000001",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "000000000",
       "000000000",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000001",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "011011100",
       "011011100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "011011100",
       "100100100",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "011100100",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011100100",
       "001001001",
       "000000000",
       "001001010",
       "000000001",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "010010010",
       "000000000",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "011011100",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011011100",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000001",
       "000001001",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "000000000",
       "001010010",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "000001001",
       "010010010",
       "000000000",
       "001001001",
       "100100101",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "100100100",
       "011011100",
       "000000000",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "100100100",
       "111111111",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "011011100",
       "011100100",
       "001001010",
       "000000000",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "011100100",
       "011100100",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "011011100",
       "011100100",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "011011100",
       "111111111",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "011100100",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "011011100",
       "100100100",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "011100100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "111111111",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "111111111",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "111111111",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "111111111",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "011100100",
       "000000000",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "000000000",
       "000000001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "011100100",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "011011100",
       "000000000",
       "000000000",
       "001010010",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "010010011",
       "000000000",
       "000000000",
       "100100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000001",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "000000001",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "010010011",
       "000000000",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "000001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "011011100",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000001",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "011011100",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "010010011",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "001010010",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "000000001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000001001",
       "000000000",
       "000000001",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "001001010",
       "010010011",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "010010011",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001001",
       "000000001",
       "000000001",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "000001001",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "100100101",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "000001001",
       "001010010",
       "001001010",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000000000",
       "000001001",
       "000000000",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "011100100",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "100100100",
       "000001001",
       "000000000",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "010010011",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "000001001",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "100100101",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001001",
       "000000000",
       "010010010",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "010010010",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "000000000",
       "001001001",
       "001001001",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "001001001",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "001001001",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "011011011",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011100",
       "100100100",
       "111111111",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "011011011",
       "011100011",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "011100011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "111111111",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "111111111",
       "011100011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "011100011",
       "111111111",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011100011",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011100011",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "011100011",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011100011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "011100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100011",
       "111111111",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "011100011",
       "011100011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100101101",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011011011",
       "011100011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100101100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001001",
       "011011011",
       "001001001",
       "001001001",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "011011011",
       "100100100",
       "100100101",
       "011011011",
       "001010010",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "001001001",
       "011011011",
       "001001001",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "100100101",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "010011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "010010010",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "010010010",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "001001001",
       "011011011",
       "010010010",
       "011011011",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001010",
       "011011011",
       "011100100",
       "100100100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100101",
       "011011100",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "100100101",
       "011011100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "010010010",
       "011011100",
       "001001001",
       "001001010",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "001010010",
       "000001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "000001001",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "010010010",
       "011100100",
       "001001010",
       "000001001",
       "010010010",
       "011011100",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001001",
       "100100101",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "100100101",
       "001001001",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "011011100",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "010010010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "010010010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "001001010",
       "010010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "001001001",
       "010010010",
       "011011100",
       "001001010",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "000001001",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "000001001",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011011",
       "001001001",
       "100100101",
       "100100100",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001001",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "100100100",
       "000001001",
       "100100101",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "100100100",
       "001010010",
       "001001001",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "010010011",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "011011100",
       "011011100",
       "001001001",
       "001001010",
       "011011100",
       "011011100",
       "001010010",
       "010010010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "000001001",
       "010010010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "100100101",
       "011011100",
       "010010010",
       "011011100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "100100100",
       "001001001",
       "011100100",
       "010010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "011100100",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "010010011",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "100100101",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "010010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "010010010",
       "000001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "010010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "010010011",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "010010011",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000001",
       "000000001",
       "000000000",
       "001001010",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000001",
       "000000000",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "000001001",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "010010011",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010011",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001010010",
       "001010010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "000001010",
       "011011100",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "100100101",
       "001001010",
       "000001010",
       "100100101",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "010010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "100100101",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001010011",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "000001010",
       "001001010",
       "100100101",
       "001001010",
       "000001001",
       "100100101",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100101",
       "001010010",
       "000001001",
       "100100101",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "000001010",
       "001001010",
       "011100101",
       "001001010",
       "000001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "010010010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "000001001",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "010010010",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "001010010",
       "011100101",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "000001010",
       "011100101",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "011100101",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "010010011",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "010010011",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "100100101",
       "001010010",
       "001001010",
       "100100101",
       "011011100",
       "001010010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "000001010",
       "001001010",
       "100100101",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "100100101",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001001",
       "010010010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "010010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001010010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000001001",
       "001010010",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "100100101",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "010010011",
       "011100100",
       "001001010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "010010011",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "000000000",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000001001",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "000001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000001",
       "000001001",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001010010",
       "011011100",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "000001001",
       "000000000",
       "000001001",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "011100100",
       "010010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "100100100",
       "011100100",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "000001001",
       "100100100",
       "001001010",
       "001001001",
       "011011100",
       "011100100",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001001",
       "100100100",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "000000001",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "001010010",
       "100100101",
       "000001001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "000000000",
       "001001010",
       "000001001",
       "010010011",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "010010011",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "010011011",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "010010011",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "000001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000001",
       "000001001",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "000001001",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "100100101",
       "001001001",
       "011011100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001010010",
       "100100100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000000000",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "010010011",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "000000001",
       "001010010",
       "001001010",
       "001010010",
       "000001001",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "100100100",
       "001010010",
       "000000000",
       "000000001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "000001001",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "000001001",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "010010010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "000001001",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001001",
       "001010010",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "000000000",
       "000000000",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010011",
       "000000001",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100101",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000001",
       "010010011",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000001",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "100100101",
       "011011011",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "000000000",
       "011100100",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "011011100",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001010011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011100",
       "011100100",
       "001001001",
       "000001001",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000001",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "000000000",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100101",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "010010011",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011011",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "010010011",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "000000000",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "010010011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "000001001",
       "001001010",
       "011100100",
       "011011100",
       "010010010",
       "011011011",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "000000001",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "010010011",
       "000000000",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "000001001",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001001",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "011100100",
       "011011100",
       "010010010",
       "011011011",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "000001001",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "000001001",
       "011100100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "000001001",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "000001001",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "010010011",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001010010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "010010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "000000000",
       "001010011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000001",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "001010011",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001001",
       "000000001",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000001010",
       "001001010",
       "000001010",
       "000000001",
       "001010010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010011",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "000000001",
       "000001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001001",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010011",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "000001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "000000000",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "010010011",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000000001",
       "000001010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001010010",
       "000000001",
       "001001010",
       "000001010",
       "010010011",
       "000001001",
       "000000001",
       "000001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "000001010",
       "001010011",
       "000001010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "000000001",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "010010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001001",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000000000",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011011",
       "001001001",
       "100100100",
       "001001010",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "000000000",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000000001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001010011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001010011",
       "000000001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "000000000",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "011100100",
       "100100100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "011011011",
       "010010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "011011100",
       "010010010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "000000000",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001001",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "001001001",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "100100100",
       "001001001",
       "000000001",
       "000001001",
       "010010011",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010011",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "000000001",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "000001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "000001001",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "000001001",
       "001010011",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "000000000",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "000000000",
       "001001010",
       "001010011",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "000001010",
       "000001010",
       "001010010",
       "000000000",
       "001001010",
       "000001010",
       "001010011",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001001",
       "000001001",
       "001010010",
       "001001010",
       "000001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "000001001",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000000000",
       "001010010",
       "000001010",
       "000001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010011",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "010010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "000001010",
       "000001010",
       "010010011",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001010010",
       "000001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "010010010",
       "011011011",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "001010010",
       "001001001",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001010011",
       "000001001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "001001001",
       "011011100",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001010011",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001010010",
       "001001001",
       "100100100",
       "001010010",
       "011100100",
       "001001001",
       "001001001",
       "011011100",
       "000000000",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001010010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "000000000",
       "011011100",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000000001",
       "001001010",
       "000001010",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "011011100",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001010010",
       "000001001",
       "001010011",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "000000000",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "010010010",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "010010011",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "000000000",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "100100101",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000000000",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100101",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "000001010",
       "000001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "000001001",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "000001001",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "011011100",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "011100100",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "100100101",
       "001001010",
       "001001010",
       "011100101",
       "000001010",
       "001001010",
       "011011100",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "000001001",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "000001001",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "010010011",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "100100101",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100101",
       "011011100",
       "011100100",
       "001001010",
       "000001001",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100101",
       "011011100",
       "011100100",
       "100100101",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "000000000",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100101",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100101",
       "011011100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100101",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100101101",
       "011011011",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011011100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "000000000",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001010010",
       "001001001",
       "011011100",
       "001010010",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "000000001",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000001",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001001",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "000001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "011011100",
       "001010010",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "000001001",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011011011",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "000001001",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001001",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001010010",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "001001001",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "011011011",
       "001001001",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "001001001",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "010010010",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "001001001",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "010010010",
       "011011011",
       "011011100",
       "001001001",
       "011011100",
       "011100100",
       "100100101",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011011100",
       "011011100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100101101",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "010011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100101101",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "000000000",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "001001010",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011011100",
       "011011100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "000000000",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "000001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100101101",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "010010010",
       "011011011",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011011011",
       "001001010",
       "011100100",
       "010010010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "011011100",
       "010010010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "010010010",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "011011100",
       "100100100",
       "100100100",
       "000001001",
       "011011100",
       "100100101",
       "001001001",
       "011011011",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011011011",
       "011100100",
       "001001010",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "001001001",
       "001001001",
       "100100101",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "100100101",
       "000001001",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001001",
       "100100101",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001010010",
       "000001001",
       "001010010",
       "001010010",
       "001010010",
       "010010010",
       "001010010",
       "000001001",
       "000000000",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "100100101",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011011011",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "010010011",
       "011100100",
       "001001010",
       "000001001",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "100100101",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "010010011",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001010010",
       "100100101",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100101",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "100100101",
       "001010010",
       "011100100",
       "000001001",
       "100100100",
       "001001001",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "011011011",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "100100101",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "100100101",
       "011011100",
       "100100101",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001010010",
       "011100100",
       "100100101",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "010010010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "100100101",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "010010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "100100101",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011100101",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "011100101",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100101",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "001010010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "100100101",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "000001001",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "010010011",
       "001001010",
       "011100100",
       "011011100",
       "010010010",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "100100101",
       "000001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001010010",
       "000001001",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000001001",
       "100100101",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "000001010",
       "001010010",
       "001001010",
       "100100101",
       "000001010",
       "011100101",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "000001010",
       "011100100",
       "001001010",
       "000001001",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010011",
       "010011100",
       "001001010",
       "010010011",
       "001001001",
       "011100100",
       "011011011",
       "010010010",
       "011100100",
       "011011011",
       "100100100",
       "000001001",
       "011011100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "000001001",
       "001010010",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "000001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "000001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "000001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011100101",
       "000001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "000001001",
       "100100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "000001001",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011100101",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "000001001",
       "011011100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "000001001",
       "001010010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "011011100",
       "001010010",
       "001001010",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "100100101",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "000001001",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "100100101",
       "001010010",
       "100100101",
       "001001001",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001001",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "010011011",
       "010010010",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "010010011",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "010010010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "010010010",
       "001001001",
       "100100101",
       "001010010",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "100100101",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "001001001",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "000001001",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "100100101",
       "001001001",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "010010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "010010011",
       "000001001",
       "001010010",
       "100100101",
       "001001010",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "100100101",
       "000001001",
       "001001010",
       "100100100",
       "000000001",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "000001001",
       "100100100",
       "001001010",
       "001001010",
       "010011011",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "010011011",
       "001010010",
       "011100100",
       "001001010",
       "000001001",
       "100100101",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100101",
       "000001001",
       "000001001",
       "100100101",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "011100100",
       "001010010",
       "100100101",
       "011100100",
       "000001001",
       "010010011",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "011100100",
       "010010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "100100101",
       "000001001",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "010010010",
       "000001001",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001001",
       "100100101",
       "010010010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "001010010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100101",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "010010010",
       "000000001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "100100101",
       "001001010",
       "000001001",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "001001010",
       "001010010",
       "011011100",
       "000001001",
       "001010010",
       "011100100",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "100100101",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "100100101",
       "000001001",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "100100101",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "100100101",
       "010010011",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "100101101",
       "001001010",
       "011011100",
       "100100101",
       "000001001",
       "011100100",
       "000001001",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "010010011",
       "011011100",
       "001001010",
       "001001010",
       "000000001",
       "100100101",
       "001001010",
       "001001010",
       "100100101",
       "001001001",
       "001010010",
       "001001001",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011011011",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "100100101",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100101",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011100",
       "000001001",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011011",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "100100101",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100101",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "000001001",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100101",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "100100101",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100101",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "000001001",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "010010010",
       "010011011",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "100100100",
       "001010010",
       "011011100",
       "001010010",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "001001001",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "000001001",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "100100100",
       "000001001",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "011011100",
       "010010010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "010010010",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "000001001",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "000001001",
       "011011100",
       "001001001",
       "100100101",
       "001001001",
       "011100100",
       "000001001",
       "100100100",
       "001001001",
       "100100101",
       "001010010",
       "001001010",
       "011011100",
       "010010010",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100101",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "000001001",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "010010011",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "100100101",
       "001001001",
       "100100101",
       "000001001",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "010010010",
       "011011100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "100100101",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100101",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "000001001",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "100100101",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "000001001",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "000001001",
       "100100100",
       "001001001",
       "011011100",
       "010010010",
       "011011100",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "000001001",
       "000000000",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011011",
       "010010010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "010010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "000001001",
       "100100101",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001010010",
       "001001010",
       "000000000",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100101",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100101",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "000001001",
       "100100101",
       "000001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "100100101",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "010010010",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "001001010",
       "000001001",
       "100100101",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "001001001",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001010010",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "100100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "011011100",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "100100100",
       "000001001",
       "100100101",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "000001001",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "010010010",
       "011100100",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011011",
       "001001001",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "001001010",
       "100100101",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "100100101",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "000001001",
       "001010010",
       "011011100",
       "011011100",
       "100100101",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "100100101",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "001001010",
       "011011100",
       "011100100",
       "100100101",
       "011011100",
       "000001001",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "000001001",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "010010010",
       "011011100",
       "001001001",
       "100100101",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "000001001",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001001",
       "011011100",
       "100100101",
       "001001001",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "010010010",
       "011011100",
       "001001001",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "001001010",
       "011011100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "000001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "011011100",
       "100100101",
       "001001001",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "000001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "100100101",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011011011",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "000001001",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011100",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "000001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "010010010",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "000001001",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100101",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "010010010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "100100101",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "001010010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "000001001",
       "100100101",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "100100100",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100101",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "100100101",
       "001001001",
       "011100100",
       "010010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "100100101",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "100100100",
       "000001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "010010010",
       "011100100",
       "011011100",
       "010010010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "001001010",
       "000001001",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "000001001",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "000001001",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100101",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "010010010",
       "011011100",
       "001010010",
       "011011100",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "011011100",
       "100100101",
       "100100100",
       "011011011",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "010010010",
       "100100100",
       "001001001",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "000001001",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "100100101",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100101",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "001010010",
       "001001010",
       "011100100",
       "100100100",
       "000000001",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "010010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001001",
       "100100101",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "001001001",
       "011011100",
       "100100100",
       "011011100",
       "001001001",
       "001010010",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011011100",
       "011011100",
       "001001001",
       "011100100",
       "011011011",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "001010010",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "010010010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "100100101",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "010010010",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "011100100",
       "001010010",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "001001010",
       "011011011",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "001001001",
       "000000000",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100101",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011011",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "011011100",
       "001010010",
       "011100100",
       "000001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "000001001",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001001010",
       "011011100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "000000000",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "010010010",
       "001001001",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "000001001",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "000001001",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "000000000",
       "011011100",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "001001010",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "010010010",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001010",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "100100101",
       "000001001",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "001001001",
       "001001001",
       "001001001",
       "011011011",
       "100100100",
       "000001001",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "000001001",
       "100100100",
       "011011011",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "000001001",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "000001001",
       "001010010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "001010010",
       "011011011",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011100100",
       "001001010",
       "001001001",
       "001001001",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "010010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "100100101",
       "011011011",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "000001001",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "100100101",
       "001001010",
       "011011100",
       "011100100",
       "010010011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "000000001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "001010010",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011011",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "000001001",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "011011011",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "000000001",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011011011",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "011011011",
       "001010010",
       "011011100",
       "011011100",
       "010010010",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011011011",
       "010010010",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "010010010",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "010010010",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001001",
       "100101101",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011011011",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "000001001",
       "011011100",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001010010",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "001010010",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "011011100",
       "001001001",
       "011011100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011011011",
       "100100100",
       "011011100",
       "001001001",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "001001001",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011011011",
       "100100100",
       "001010010",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "001010010",
       "000001001",
       "011011011",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011011100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "001010001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "000001001",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001010010",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "000001001",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "010010010",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "000001001",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011100011",
       "001010010",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "001001001",
       "011011011",
       "100100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "010010010",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100101101",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "000001001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001010001",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010001",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "000001001",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001001001",
       "001001010",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "010010010",
       "011011011",
       "000001001",
       "011100100",
       "001010010",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "010010010",
       "011011011",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "000001001",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "000001001",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "010010010",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "011011011",
       "100101101",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "010010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001010001",
       "011100011",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "010010010",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "001010010",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "010010010",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "000001001",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "010010010",
       "011011011",
       "011100100",
       "011100100",
       "000000000",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100011",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "010011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001001",
       "001010010",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001010010",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001010010",
       "011011100",
       "011011011",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "011011011",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "010010011",
       "001001001",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "000001001",
       "010010010",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "010010010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "010010010",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001001001",
       "010010010",
       "000001001",
       "001001001",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "000001001",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "001010010",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "001010010",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "001001001",
       "010010010",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100101101",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "010010010",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "010010010",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "010010010",
       "001001001",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100101101",
       "011011011",
       "011011100",
       "011011100",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001010",
       "000001001",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100101",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "001001001",
       "001001001",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "010010010",
       "010011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "001001001",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100101",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "001001001",
       "100100100",
       "111111111",
       "011100100",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "001001001",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "001001001",
       "001001001",
       "011100100",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "001010001",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001001",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001010010",
       "001001001",
       "011011011",
       "100100101",
       "011011011",
       "000001001",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "010010010",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "010010010",
       "001001001",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "001010001",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100101",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "001010001",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100101",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "000001001",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "000001001",
       "001010010",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "010010010",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "111111111",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "011100011",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011011011",
       "001001010",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011011100",
       "001010010",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "010010010",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100101",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "010010010",
       "011011100",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "001001001",
       "001001001",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "001001001",
       "001001001",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "010010010",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "010010010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "011011100",
       "111111111",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "000001001",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011011100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001010010",
       "000001001",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "001010010",
       "001010010",
       "011100100",
       "001010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100101",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "001010010",
       "011011011",
       "001010010",
       "011011100",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "100100101",
       "011011100",
       "001001001",
       "010010010",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "001010010",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "010010010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "010010010",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100101",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011011011",
       "001001001",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001001001",
       "010010010",
       "000001001",
       "001001010",
       "001001001",
       "000001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "010010010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "000000000",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "000000000",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "001001001",
       "000000000",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "001001001",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "010010010",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "010010010",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100101",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "010010010",
       "011100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "011011100",
       "001001010",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001001001",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "010010010",
       "011011100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "011011100",
       "001001010",
       "100100100",
       "011011011",
       "010010010",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "001001010",
       "011011011",
       "100100101",
       "011011011",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100101",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "001001001",
       "100100101",
       "011011100",
       "001010010",
       "011011011",
       "011100100",
       "001010010",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "010010010",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011011011",
       "010010010",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011011011",
       "001010010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011011",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "011011011",
       "010010010",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "100100100",
       "011011011",
       "100100100",
       "000001001",
       "100100100",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "001010010",
       "011100100",
       "011100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011011100",
       "001010010",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011011100",
       "011011100",
       "001001001",
       "100100101",
       "011011100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "011011100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "100100100",
       "000001001",
       "011100100",
       "100100100",
       "011011100",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "000001001",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "011011100",
       "001010010",
       "000001001",
       "100100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "000001001",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "011011011",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011011100",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001010010",
       "001001001",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "001010010",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001001010",
       "011100100",
       "011100100",
       "010010010",
       "010011011",
       "100100100",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "001010010",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "011011011",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "011011100",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "100100100",
       "000001001",
       "001001010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "100100100",
       "001001001",
       "011011100",
       "100100100",
       "001001001",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "100100100",
       "001001001",
       "001001010",
       "100100100",
       "011011100",
       "001001010",
       "011100100",
       "011011100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "000001001",
       "011100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "010010010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "000001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "010010010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000001001",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "011100100",
       "001001001",
       "001010010",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "011100100",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001001010",
       "100100100",
       "001010010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "001010010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "000001001",
       "001001001",
       "001010010",
       "011011100",
       "011011100",
       "010010010",
       "011100100",
       "001010010",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011011011",
       "001001010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001010010",
       "001001010",
       "011100100",
       "010010010",
       "100100100",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "001001001",
       "001001001",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011011100",
       "001001001",
       "011100100",
       "001010010",
       "011100100",
       "001001001",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "100100100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001001",
       "011100100",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001001",
       "001010010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011100",
       "011011100",
       "001010010",
       "011100100",
       "000001001",
       "011100100",
       "001001010",
       "011011100",
       "010010010",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001010010",
       "011100100",
       "001001010",
       "001001001",
       "001010010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "011100100",
       "001010010",
       "011011011",
       "010010010",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "011100100",
       "001010010",
       "011011100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001001",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "100100100",
       "001001001",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "011100100",
       "001001001",
       "001010010",
       "100100100",
       "001001010",
       "001001001",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011100",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011100",
       "011011011",
       "100100100",
       "111111111",
       "011011100",
       "011100100",
       "111111111",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "011011100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "011011100",
       "011011100",
       "011100100",
       "100100101",
       "011011100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "011011100",
       "111111111",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100101",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "111111111",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "100100101",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "111111111",
       "011100100",
       "011011100",
       "011011100",
       "111111111",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "011011100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "011011100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100101",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "011011100",
       "111111111",
       "011100100",
       "011011011",
       "011011100",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011100",
       "111111111",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011100011",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "111111111",
       "011011100",
       "100100100",
       "011011011",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "100100011",
       "100100011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100011",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "011011100",
       "111111111",
       "011011100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011100100",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011011011",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011100011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "111111111",
       "011011011",
       "011100011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "011100100",
       "011100011",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "111111111",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "011100011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100011",
       "011011011",
       "011100100",
       "011100011",
       "011100011",
       "111111111",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011100011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011011011",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100011",
       "100100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "011100100",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "011100011",
       "111111111",
       "011100011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100011",
       "011100100",
       "011100011",
       "011011011",
       "111111111",
       "011100011",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011100011",
       "100100100",
       "011100011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100011",
       "100100100",
       "011100011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "111111111",
       "011100100",
       "011100011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011100011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "001001001",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011100100",
       "111111111",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011011011",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001001010",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "001001001",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100101",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "001010010",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011011011",
       "001010010",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "001001001",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "111111111",
       "100100100",
       "111111111",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "001001001",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001001",
       "011011100",
       "011100100",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "001001001",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "111111111",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "001001010",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011011",
       "001001001",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "011011011",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "011011011",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "011011100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001001001",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "001001010",
       "011100100",
       "011011100",
       "011100100",
       "011011100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "100100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "001010010",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011011100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100101",
       "011011011",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "001001001",
       "011100100",
       "011100100",
       "011011100",
       "011100100",
       "011011011",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "100100100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "100100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "001010010",
       "100100100",
       "011011100",
       "100100100",
       "100100100",
       "011011100",
       "100100100",
       "011011011",
       "100100101",
       "011011011",
       "100100100",
       "011100100",
       "011011011",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "100100100",
       "100100100",
       "011011011",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "100100101",
       "011011100",
       "011100100",
       "100100100",
       "011011100",
       "011011100",
       "011100100",
       "100100100",
       "011011011",
       "011011100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011011100",
       "001001001",
       "011011100",
       "100100100",
       "011011100",
       "011100100",
       "011100100",
       "100100100",
       "011011100",
       "011100100",
       "011011100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "100100100",
       "011100100",
       "100100100",
       "011100100",
       "011100100",
       "011100100",
       "011100100",
       "011011100",
       "100100100",
       "011011100",
       "011011011",
       "100100100",
       "011100100",
       "100100100",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "111111111",
       "011011100",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001010010",
       "000000000",
       "111111111",
       "011100100",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "010010011",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "011100100",
       "111111111",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "010010010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "111111111",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "111111111",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "011011100",
       "100100100",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "011011100",
       "100100100",
       "001001010",
       "001010010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "111111111",
       "010010010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "010010011",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "011011100",
       "011011100",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "111111111",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "010010011",
       "011100100",
       "001001010",
       "000000000",
       "000001001",
       "001010010",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "100100100",
       "100100100",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "100100100",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "010010011",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "100100101",
       "000000000",
       "000000000",
       "000001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000001001",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "010010010",
       "000001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000001001",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "000000001",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000001001",
       "001010010",
       "000000000",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "010010011",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "001001001",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000001",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "000001001",
       "000000001",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "100100101",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "000000000",
       "100100100",
       "011011100",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001010",
       "001010010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "010010010",
       "001001001",
       "000000000",
       "010010010",
       "001001001",
       "001001010",
       "001001010",
       "000000000",
       "100100100",
       "011100100",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "001001001",
       "010010010",
       "000000000",
       "010010010",
       "001001010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "011011100",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "010010010",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "011011100",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "111111111",
       "001010010",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "011100100",
       "010010010",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001001010",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "100100100",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "001001010",
       "000000001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "010010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "011100100",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "010010010",
       "010010010",
       "000001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "010010010",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "011100100",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "001001010",
       "001010010",
       "001010010",
       "001001001",
       "001001010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001001",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "001001001",
       "001001001",
       "001001010",
       "011011100",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "000000001",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "010010010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "001001010",
       "001001001",
       "001001010",
       "001001010",
       "001001010",
       "000001001",
       "001001010",
       "001010010",
       "001001001",
       "001001010",
       "001010010",
       "000001001",
       "001010010",
       "001001010",
       "001001001",
       "001010010",
       "001010010",
       "001001001",
       "001001001",
       "001010010",
       "001001001",
       "100100100",
       "000000000",
       "001001010",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "010010010",
       "001001001",
       "001001001",
       "010010010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "011100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "100100100",
       "001001001",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "010010010",
       "011011100",
       "001001010",
       "001001001",
       "100100100",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "011011100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "010010010",
       "011100100",
       "001001001",
       "001001010",
       "001001001",
       "011100100",
       "001001001",
       "100100100",
       "001001001",
       "001001001",
       "001010010",
       "100100100",
       "001001010",
       "010010010",
       "011100100",
       "001001001",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "100100100",
       "001001001",
       "001001001",
       "100100100",
       "001001010",
       "010010010",
       "011011100",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011100",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "001001010",
       "100100100",
       "001001010",
       "011011100",
       "010010010",
       "001001001",
       "011100100",
       "001001001",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001001",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "100100100",
       "001010010",
       "001001001",
       "001001010",
       "011100100",
       "001001001",
       "001001010",
       "011011100",
       "001001010",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001001010",
       "011100100",
       "001001010",
       "001010010",
       "001001001",
       "100100101",
       "001001001",
       "001001001",
       "011100100",
       "001001010",
       "001001010",
       "011100100",
       "001001010",
       "000000001",
       "001010010",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000001",
       "001001001",
       "100100100",
       "001001001",
       "001001001",
       "001001001",
       "100100100",
       "000001001",
       "001001010",
       "100100101",
       "001001001",
       "011011100",
       "001001010",
       "001001010",
       "001001010",
       "011011100",
       "001010010",
       "011100100",
       "001001001",
       "001010010",
       "001001001",
       "001010010",
       "100100100",
       "001001001",
       "001001010",
       "011100100",
       "001010010",
       "001001001",
       "100100100",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "011011100",
       "001001001",
       "100100100",
       "001001010",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001010001",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000001",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001010010",
       "001001001",
       "000000000",
       "000000000",
       "010010010",
       "001001001",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "001001001",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001010001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000001",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "001001010",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "010010010",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "010010010",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "010010010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001010010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "001001010",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "001001001",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

