------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : mapadeverdadpeque.ppm 
--- Filas    : 256 
--- Columnas : 256 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_mapadeverdadpeque is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(16-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_mapadeverdadpeque;


architecture BEHAVIORAL of ROM_RGB_9b_mapadeverdadpeque is
  signal addr_int  : natural range 0 to 2**16-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "111111111",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "001001010",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "001010010",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "001001010",
       "011011011",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "001010010",
       "011011011",
       "001001010",
       "001010010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001010010",
       "100100100",
       "001010010",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "011011011",
       "001010010",
       "011011011",
       "001010010",
       "001001010",
       "100100100",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001010010",
       "100100100",
       "001001010",
       "001001010",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "001010010",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "111111111",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "111111111",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "001001010",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "111111111",
       "100100100",
       "111111111",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "001001010",
       "100100100",
       "001010010",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "111111111",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "001010010",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "001001010",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "100100100",
       "100100100",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "001001010",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "011011011",
       "100100100",
       "011011011",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "111111111",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "100100100",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "011011011",
       "001001010",
       "011011011",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001010010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010",
       "001001010"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

