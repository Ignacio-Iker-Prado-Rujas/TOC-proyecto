--------------------------------------------------------------------------------
-- Felipe Machado Sanchez
-- Departameto de Tecnologia Electronica
-- Universidad Rey Juan Carlos
-- http://gtebim.es/~fmachado
--

------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    Clk  :  senal de reloj
--    Addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    Dout : dato de 3 bits, indica el tipo de pared:
--
--        "000": pared interior o pasillo  (no se pinta)
--        "001": pared vertical                    |
--        "010": pared horizontal                  _
--                                                 _ 
--        "011": esquina superior izquierda       |
--        "100": esquina inferior izquierda       |_
--                                                 _ 
--        "101": esquina superior derecha           |
--        "110": esquina inferior derecha          _|
--

--  Esta ROM idica el tipo de esquina, esto se saca a partir de las paredes
--  del laberinto, laberinto de 32 columnas x 30 filas, pero como la mitad
--  derecha es sim�trica con la izquierda, no es necesario repetirla
--  por lo tanto tiene 16 columnas x 30 filas = 480 elementos


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;

library WORK;
use WORK.PACMAN_PKG.ALL;

entity ROM_paredlaberin is
  port (
    clk   : in  std_logic;   
    addr : in  std_logic_vector(c_nb_cuad_num-2 downto 0);
    dout : out std_logic_vector(2 downto 0)
  );
end ROM_paredlaberin;

architecture BEHAVIORAL of ROM_paredlaberin is
  type memostruct is array (natural range<>) of
                   std_logic_vector(2 downto 0);

  constant img : memostruct := (
 -- F     E     D     C     B     A     9     8     7     6     5     4     3     2     1     0
  "011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101", -- 0
  "001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001", -- 1
  "001","000","011","010","010","101","000","011","010","010","010","010","010","101","000","001", -- 2
  "001","000","001","000","000","001","000","001","000","000","000","000","000","001","000","001", -- 3
  "001","000","100","010","010","110","000","100","010","010","010","010","010","110","000","100", -- 4
  "001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000", -- 5
  "001","000","011","010","010","101","000","011","101","000","011","010","010","010","010","010", -- 6
  "001","000","100","010","010","110","000","001","001","000","100","010","010","010","010","101", -- 7
  "001","000","000","000","000","000","000","001","001","000","000","000","000","000","000","001", -- 8
  "100","010","010","010","010","101","000","001","100","010","010","010","010","101","000","001", -- 9
  "000","000","000","000","000","001","000","001","011","010","010","010","010","110","000","100", --10
  "000","000","000","000","000","001","000","001","001","000","000","000","000","000","000","000", --11
  "010","010","010","010","010","110","000","100","110","000","011","010","010","010","000","000", --12
  "000","000","000","000","000","000","000","000","000","000","001","000","000","000","000","000", --13
  "010","010","010","010","010","101","000","011","101","000","001","000","000","000","000","000", --14
  "000","000","000","000","000","001","000","001","001","000","100","010","010","010","010","010", --15
  "000","000","000","000","000","001","000","001","001","000","000","000","000","000","000","000", --16
  "000","000","000","000","000","001","000","001","001","000","011","010","010","010","010","010", --17
  "011","010","010","010","010","110","000","100","110","000","100","010","010","010","010","101", --18
  "001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001", --19
  "001","000","011","010","010","101","000","011","010","010","010","010","010","101","000","001", --20
  "001","000","100","010","101","001","000","100","010","010","010","010","010","110","000","100", --21 
  "001","000","000","000","001","001","000","000","000","000","000","000","000","000","000","000", --22
  "100","010","101","000","001","001","000","011","101","000","011","010","010","010","010","010", --23
  "011","010","110","000","100","110","000","001","001","000","100","010","010","010","010","101", --24
  "001","000","000","000","000","000","000","001","001","000","000","000","000","000","000","001", --25
  "001","000","011","010","010","010","010","110","100","010","010","010","010","101","000","001", --26
  "001","000","100","010","010","010","010","010","010","010","010","010","010","110","000","100", --27
  "001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000", --28
  "100","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"  --29

    );

begin

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= img(to_integer(unsigned(addr)));
    end if;
  end process;

end BEHAVIORAL;

