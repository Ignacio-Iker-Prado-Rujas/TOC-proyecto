------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : lab.ppm 
--- Filas    : 256 
--- Columnas : 128 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_lab is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(15-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_lab;


architecture BEHAVIORAL of ROM_RGB_9b_lab is
--  signal addr_int  : natural range 0 to 2**15-1;
--  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
--  constant filaimg : memostruct := (
--     --"RRRGGGBBB"
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "111111111",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "111111111",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "100100100",
--       "100100100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100",
--       "000000100"
--        );

begin

  --addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      --dout <= filaimg(addr_int);
		dout <= "000000100";
    end if;
  end process;

end BEHAVIORAL;

