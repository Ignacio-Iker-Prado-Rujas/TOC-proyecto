--------------------------------------------------------------------------------
-- Felipe Machado Sanchez
-- Departameto de Tecnologia Electronica
-- Universidad Rey Juan Carlos
-- http://gtebim.es/~fmachado
--
------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 1 bit de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;

library WORK;
use WORK.PINTAROM_PKG.ALL;

entity ROM1b_16x16 is
  port (
    clk  : in  std_logic;  
    addr : in  std_logic_vector(7 downto 0);
    dout : out std_logic 
  );
end ROM1b_16x16;


architecture BEHAVIORAL of ROM1b_16x16 is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic;

  constant img : memostruct := (
 -- 0   1   2   3   4   5   6   7   8   9  10  11  12  13  14  15
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 0
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 1
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 2
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 3
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 4
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 5
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 6
   '1','0','1','0','1','0','1','0','1','0','1','0','1','0','1','0', -- 7
   '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1', -- 8
   '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', -- 9
   '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1', --10
   '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', --11
   '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1', --12
   '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', --13
   '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1', --14
   '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'  --15
  );

begin

  Addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= img(addr_int);
    end if;
  end process;

end BEHAVIORAL;

