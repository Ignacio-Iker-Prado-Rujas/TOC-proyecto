------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : patron_100x100_gris.pgm 
--- Filas    : 100 
--- Columnas : 100 
--- Color    :  8 bits



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM8b_patron_100x100_gris is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(14-1 downto 0);
    dout : out std_logic_vector(8-1 downto 0) 
  );
end ROM8b_patron_100x100_gris;


architecture BEHAVIORAL of ROM8b_patron_100x100_gris is
  signal addr_int  : natural range 0 to 2**14-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
       "10110110",
       "11111111",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "01101010",
       "11111111",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "10110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11101000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110000",
       "01110000",
       "01110000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "01100110",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "10100100",
       "11111111",
       "10100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "00000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

