------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : Joyride.ppm 
--- Filas    : 64 
--- Columnas : 32 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_Joyride is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(11-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_Joyride;


architecture BEHAVIORAL of ROM_RGB_9b_Joyride is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111110110",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111101110",
       "111110110",
       "100010010",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011010001",
       "100011001",
       "100010001",
       "100011010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111110110",
       "110101101",
       "011010010",
       "111110110",
       "111110110",
       "010001001",
       "101011011",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "110101101",
       "100011010",
       "011010001",
       "100011001",
       "101100010",
       "100010001",
       "101011011",
       "110100100",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "110101101",
       "100011011",
       "100011011",
       "100011011",
       "010001001",
       "101011011",
       "100011010",
       "011010010",
       "100010010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110111",
       "100011011",
       "010001000",
       "101101011",
       "111110011",
       "111110011",
       "101100001",
       "100011001",
       "100010010",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "100010011",
       "010001000",
       "010001000",
       "010001001",
       "100011010",
       "010001000",
       "010001000",
       "101011011",
       "100010010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "001000000",
       "100011001",
       "101100010",
       "111110010",
       "111101001",
       "111110010",
       "111110100",
       "010001000",
       "111101101",
       "111110110",
       "110101101",
       "111101101",
       "001000000",
       "100010010",
       "011010010",
       "011010010",
       "100011011",
       "011010001",
       "100010010",
       "101011011",
       "100010010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011001001",
       "101011011",
       "101100010",
       "011011000",
       "110100001",
       "101100000",
       "110101001",
       "111111011",
       "010001000",
       "111110101",
       "111111110",
       "001000000",
       "010001000",
       "011010010",
       "011010010",
       "011010010",
       "011010001",
       "100011010",
       "100010010",
       "100010010",
       "100010010",
       "011010010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "010000000",
       "101100011",
       "010001000",
       "100100001",
       "110101001",
       "110101000",
       "101100000",
       "111110011",
       "011010001",
       "001000000",
       "010001000",
       "100011011",
       "011010010",
       "100010010",
       "011010001",
       "011010001",
       "010001000",
       "010001000",
       "010001000",
       "010001001",
       "010000000",
       "011001010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110111",
       "010001001",
       "110100100",
       "011010001",
       "001000000",
       "101100001",
       "110101000",
       "110100000",
       "110101000",
       "110101001",
       "011010000",
       "011010001",
       "011010010",
       "100011010",
       "011010001",
       "011010010",
       "010001001",
       "010001000",
       "010000000",
       "010001000",
       "010000000",
       "010001001",
       "010001001",
       "010000001",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "110100100",
       "010001001",
       "110101100",
       "011001000",
       "101100010",
       "100011000",
       "110101000",
       "110101000",
       "110100000",
       "110101001",
       "011010000",
       "010001000",
       "100010010",
       "011010001",
       "011001001",
       "011001001",
       "010001000",
       "010001000",
       "001000000",
       "001000000",
       "001000000",
       "001000000",
       "001000000",
       "101011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "100010010",
       "100011011",
       "100010010",
       "101011011",
       "111110101",
       "100011000",
       "110101001",
       "110101000",
       "110101000",
       "110101001",
       "011010000",
       "001000000",
       "011010001",
       "011010001",
       "011001001",
       "010001000",
       "010001000",
       "010001000",
       "010000000",
       "010001000",
       "010000000",
       "010000000",
       "001000000",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101011010",
       "110100100",
       "011001001",
       "111110110",
       "111110100",
       "100011000",
       "110101001",
       "110101000",
       "110101000",
       "110101001",
       "011010000",
       "001000000",
       "010001001",
       "011010001",
       "010001000",
       "010001000",
       "010001000",
       "001000000",
       "100011010",
       "101011011",
       "100011010",
       "100010010",
       "010000000",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101011011",
       "101011011",
       "110101101",
       "111110110",
       "111110101",
       "011010000",
       "100100001",
       "100100000",
       "101100000",
       "101100001",
       "010001000",
       "001000000",
       "011010001",
       "011001001",
       "010001000",
       "010001000",
       "010001000",
       "001000000",
       "111110101",
       "111111110",
       "111110101",
       "111110101",
       "011010010",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "011001001",
       "100010010",
       "101011011",
       "111110110",
       "111110110",
       "001000000",
       "011010000",
       "010010000",
       "100011000",
       "100011000",
       "001000000",
       "010000000",
       "011010001",
       "010001000",
       "010001000",
       "010001000",
       "010001000",
       "010001000",
       "111110110",
       "111111110",
       "111110101",
       "111110101",
       "101011011",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "100011010",
       "101011010",
       "111101110",
       "111101110",
       "111101101",
       "100011010",
       "110101011",
       "001000000",
       "101100010",
       "111110100",
       "001000000",
       "001000000",
       "010001000",
       "010001000",
       "010001000",
       "010001000",
       "010000000",
       "011001001",
       "111110101",
       "011010001",
       "011010001",
       "101011010",
       "100010010",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "100010010",
       "100010010",
       "111110110",
       "111101110",
       "111101101",
       "010001000",
       "111111101",
       "100011001",
       "011010000",
       "100011010",
       "001000000",
       "010001000",
       "010001000",
       "010001000",
       "010001000",
       "010001000",
       "010000000",
       "011001001",
       "111110101",
       "100011001",
       "011010001",
       "011001001",
       "011001001",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101011100",
       "100010010",
       "101011011",
       "111101110",
       "111101110",
       "111110110",
       "011010001",
       "101101011",
       "100100010",
       "001001000",
       "010010001",
       "001000000",
       "010001000",
       "010001000",
       "010001000",
       "010001001",
       "010001001",
       "010000000",
       "010001000",
       "111110101",
       "110100011",
       "011010001",
       "011001001",
       "011001001",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011010010",
       "100010010",
       "111101101",
       "111101101",
       "111101101",
       "111110110",
       "100011011",
       "010001000",
       "011010001",
       "010010001",
       "100011011",
       "001000000",
       "010001000",
       "010001001",
       "010001000",
       "010001001",
       "010001001",
       "010000000",
       "011010001",
       "111110101",
       "101100011",
       "011010001",
       "011010001",
       "011001001",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110101",
       "101011011",
       "100010010",
       "111101101",
       "111101110",
       "111101101",
       "111110110",
       "100011011",
       "000000000",
       "000000000",
       "100100100",
       "110110101",
       "010001001",
       "001000000",
       "010001000",
       "010001000",
       "010000000",
       "010001000",
       "001000000",
       "101100011",
       "111101100",
       "100010001",
       "010001000",
       "010001001",
       "100010010",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110101",
       "101011011",
       "011001001",
       "111101101",
       "111101110",
       "111101110",
       "111110110",
       "100010011",
       "010001001",
       "010010001",
       "110110110",
       "111111110",
       "100100011",
       "001000000",
       "011001001",
       "010000000",
       "001000000",
       "010000000",
       "001000000",
       "111110101",
       "100011010",
       "100011010",
       "110101101",
       "000000000",
       "011001001",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "100011011",
       "101011011",
       "111101101",
       "111101101",
       "111101110",
       "111101110",
       "111110111",
       "001001001",
       "011011011",
       "111111110",
       "111111110",
       "101100100",
       "001000000",
       "010001001",
       "010000000",
       "111110110",
       "010001000",
       "001000000",
       "111110101",
       "110101100",
       "110101100",
       "111110110",
       "001000000",
       "011001010",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "100010010",
       "100010010",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111110111",
       "001000000",
       "101100100",
       "101100100",
       "011011010",
       "101101100",
       "001000000",
       "001000000",
       "100011011",
       "111110110",
       "100011010",
       "011001000",
       "111110101",
       "111110101",
       "110110101",
       "111110110",
       "000000000",
       "101011011",
       "101011011",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "100010010",
       "101011010",
       "101011011",
       "111110110",
       "111101110",
       "111101110",
       "111110111",
       "010001001",
       "101101100",
       "100011011",
       "011010010",
       "101100100",
       "010010001",
       "001000000",
       "111101101",
       "101100011",
       "101100011",
       "100011010",
       "111110101",
       "111111110",
       "111110101",
       "111110110",
       "010001001",
       "110101101",
       "100010010",
       "111100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011001001",
       "101011011",
       "011010001",
       "111101101",
       "111110110",
       "111110110",
       "101100100",
       "011010010",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "011010010",
       "001000000",
       "111110110",
       "101100011",
       "101100011",
       "101011010",
       "111101100",
       "111111110",
       "111110101",
       "111110110",
       "100100011",
       "111110101",
       "101011011",
       "110011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "101011010",
       "100011010",
       "100011010",
       "110101101",
       "110101101",
       "001000000",
       "010010001",
       "100011011",
       "110101101",
       "110110101",
       "101101100",
       "100011010",
       "001000000",
       "111110101",
       "111110101",
       "101011010",
       "100011010",
       "110101100",
       "111110101",
       "111111110",
       "111110110",
       "111110101",
       "111110101",
       "101011011",
       "101011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011001001",
       "011001000",
       "110100011",
       "011001000",
       "010001000",
       "010001000",
       "001001000",
       "010010001",
       "010010010",
       "101101100",
       "100100011",
       "100100011",
       "100011011",
       "001000000",
       "101100100",
       "111111110",
       "110101100",
       "100011010",
       "100011010",
       "111110101",
       "111111110",
       "101100100",
       "101100100",
       "101100011",
       "011001001",
       "110100100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011001001",
       "010000000",
       "111101100",
       "110101011",
       "111110101",
       "011010001",
       "010001000",
       "110101101",
       "011011010",
       "101101100",
       "011011010",
       "001001001",
       "001001001",
       "000000000",
       "010001001",
       "110101101",
       "111111110",
       "100011011",
       "100011010",
       "110101100",
       "110101100",
       "101100011",
       "011010001",
       "101100011",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "010001000",
       "101100011",
       "101011010",
       "111101100",
       "011010001",
       "001000000",
       "100100011",
       "011011011",
       "101101100",
       "011011010",
       "101100100",
       "010010001",
       "000000000",
       "001000000",
       "010010010",
       "011011011",
       "011010010",
       "100011011",
       "101100100",
       "110100100",
       "101100011",
       "011010001",
       "101100100",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101100100",
       "010000000",
       "101100011",
       "011010001",
       "110100011",
       "010001000",
       "010001000",
       "011011010",
       "011011011",
       "101101100",
       "011011010",
       "101100100",
       "010010001",
       "001001001",
       "001001001",
       "010001001",
       "010001001",
       "010001001",
       "011010010",
       "101100011",
       "101100100",
       "101100011",
       "011010010",
       "100011011",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "001000000",
       "101011011",
       "011010001",
       "101100011",
       "010001000",
       "010001000",
       "011010010",
       "011011011",
       "101101100",
       "100011011",
       "100011011",
       "001001001",
       "001001001",
       "010001001",
       "010010010",
       "011010010",
       "010001001",
       "010001001",
       "100011011",
       "100011011",
       "100011011",
       "011001001",
       "110100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "010000000",
       "011010010",
       "010001001",
       "011010010",
       "010001000",
       "010001000",
       "011010010",
       "100011011",
       "101100100",
       "011011010",
       "010010010",
       "001001001",
       "001000001",
       "010001010",
       "011010011",
       "101100101",
       "011010010",
       "010001001",
       "011010010",
       "001000001",
       "011010010",
       "011010010",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "101011100",
       "010000000",
       "010000000",
       "010001000",
       "001000000",
       "001001000",
       "011011010",
       "011011010",
       "101101100",
       "011011010",
       "011011010",
       "001001001",
       "001000001",
       "010001010",
       "100011011",
       "111111110",
       "100011011",
       "010001001",
       "100011011",
       "001000000",
       "011011011",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111110110",
       "111110111",
       "010001001",
       "000000000",
       "101100011",
       "100011001",
       "101101011",
       "100011010",
       "010010001",
       "001001000",
       "001001001",
       "010001010",
       "101101100",
       "111111110",
       "110101100",
       "100011011",
       "110101100",
       "100011010",
       "010001001",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "000000000",
       "011010001",
       "111110100",
       "100100001",
       "010010000",
       "100100010",
       "001001000",
       "010001010",
       "001001001",
       "101100100",
       "111111110",
       "111111110",
       "101100011",
       "011010010",
       "101100011",
       "110101100",
       "010001001",
       "101011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "010001000",
       "010010000",
       "111110011",
       "110101010",
       "010001000",
       "011011001",
       "010010000",
       "011010010",
       "001001001",
       "011010001",
       "111110101",
       "111110101",
       "111101100",
       "101100011",
       "110101100",
       "111111110",
       "100011010",
       "101011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "010010001",
       "010001000",
       "100100001",
       "111110100",
       "100011000",
       "010010000",
       "010010000",
       "010010001",
       "010010001",
       "010001000",
       "110101100",
       "111101100",
       "111110101",
       "111110101",
       "111110101",
       "111111101",
       "110101100",
       "101011011",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010001001",
       "010001001",
       "001001000",
       "010001000",
       "110110100",
       "101101010",
       "010001000",
       "010001000",
       "001001000",
       "011010010",
       "010010001",
       "011010010",
       "101100011",
       "111110101",
       "111110101",
       "111110101",
       "111110101",
       "110101100",
       "101011011",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "010010001",
       "001000000",
       "001000000",
       "001001000",
       "011011001",
       "101101011",
       "010010000",
       "001001000",
       "000000000",
       "010010010",
       "011010010",
       "001001001",
       "011010010",
       "110100100",
       "110101101",
       "110100100",
       "110100100",
       "101011011",
       "101011100",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110111",
       "100011011",
       "001000000",
       "000000000",
       "000000000",
       "001000000",
       "000000000",
       "000000000",
       "001001001",
       "001001001",
       "001001001",
       "001000001",
       "001000000",
       "100010011",
       "100011011",
       "100010010",
       "011010010",
       "011001001",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "100011100",
       "010001001",
       "001001001",
       "010010001",
       "000000000",
       "010010001",
       "000000000",
       "010001010",
       "010010010",
       "001001010",
       "001001001",
       "001000001",
       "010001010",
       "001000000",
       "110100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "100011100",
       "010001001",
       "010010001",
       "100011011",
       "001000000",
       "010010010",
       "010010010",
       "011011011",
       "001000001",
       "001001001",
       "001001001",
       "001001010",
       "001001001",
       "000000000",
       "110100101",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101011100",
       "010001001",
       "010010001",
       "100011011",
       "001001000",
       "010010010",
       "010010010",
       "110110110",
       "011011011",
       "000000001",
       "001001010",
       "010010011",
       "001001010",
       "000000000",
       "110100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "101011100",
       "010001001",
       "010010001",
       "100011011",
       "001001000",
       "010010001",
       "010001001",
       "111111111",
       "101101101",
       "000000001",
       "010010011",
       "010010011",
       "010001010",
       "000000000",
       "101100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "100011011",
       "010001001",
       "010010001",
       "011011011",
       "001001000",
       "010010001",
       "001001001",
       "111110111",
       "101100101",
       "001000001",
       "010010011",
       "010010011",
       "010001010",
       "000000000",
       "101100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "001000000",
       "010001001",
       "010001001",
       "010010010",
       "001001000",
       "010001001",
       "001001001",
       "111110111",
       "101100101",
       "000000001",
       "011011100",
       "010010011",
       "001001010",
       "000000000",
       "101100101",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "001001001",
       "011011011",
       "001001000",
       "010010001",
       "001000000",
       "000000000",
       "001001001",
       "111111111",
       "101100101",
       "000000001",
       "010010011",
       "010010011",
       "000000000",
       "011010011",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "001000000",
       "011010010",
       "011011011",
       "011011011",
       "010010010",
       "010010001",
       "001000000",
       "100011100",
       "101101101",
       "001000001",
       "011011011",
       "010010011",
       "000000000",
       "010010010",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011010010",
       "001000000",
       "100100011",
       "100100011",
       "011011010",
       "010010010",
       "001001001",
       "110101110",
       "110100101",
       "000000001",
       "010010011",
       "001001010",
       "000000000",
       "010010010",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "110101101",
       "001000000",
       "010010010",
       "010010010",
       "010001001",
       "001001001",
       "100011011",
       "111110111",
       "110101110",
       "100011100",
       "001001001",
       "000000000",
       "000000000",
       "010001010",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "011010010",
       "011010010",
       "001000000",
       "001000000",
       "001001001",
       "111110110",
       "111101110",
       "111101110",
       "111110111",
       "001001001",
       "000000000",
       "000000000",
       "001000001",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111110111",
       "001000001",
       "001000001",
       "101011100",
       "111110110",
       "111101110",
       "111101110",
       "111110110",
       "101100100",
       "000000000",
       "000000000",
       "010001001",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "111110110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111111111",
       "000000000",
       "000000000",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111110110",
       "110101101",
       "010001010",
       "111110111",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "110100101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101101",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110",
       "111101110"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

