------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : jetpack-joyride-16x32-aire.ppm 
--- Filas    : 32 
--- Columnas : 16 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_Joyride is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(9-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_Joyride;


architecture BEHAVIORAL of ROM_RGB_9b_Joyride is
  signal addr_int  : natural range 0 to 2**9-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "100100010",
       "100100001",
       "111111110",
       "111111111",
       "111111111",
       "011010001",
       "011001001",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010001000",
       "011010000",
       "111111100",
       "100100001",
       "100100001",
       "111111110",
       "001000000",
       "011010001",
       "011001001",
       "011001001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010000000",
       "011001000",
       "101011000",
       "111110010",
       "101101010",
       "101101010",
       "011010001",
       "011010001",
       "011010001",
       "011010010",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "100010000",
       "101011000",
       "110101001",
       "110101010",
       "001000000",
       "100011010",
       "011010001",
       "001000000",
       "001000000",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "101011001",
       "110101010",
       "110100001",
       "101100010",
       "001000000",
       "011010001",
       "010000000",
       "010001000",
       "011010001",
       "100011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010001000",
       "011001000",
       "011001000",
       "100010000",
       "100011000",
       "101011010",
       "001000000",
       "010001001",
       "001000000",
       "110100100",
       "111111110",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001001000",
       "010001000",
       "111111110",
       "100011001",
       "100011001",
       "100011001",
       "001000000",
       "010001000",
       "001000000",
       "111101101",
       "100010010",
       "100010010",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011010",
       "010001000",
       "111111110",
       "011010001",
       "011010001",
       "010001001",
       "001000000",
       "010001001",
       "001000000",
       "111110101",
       "010001000",
       "011001001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001001000",
       "001000000",
       "111111111",
       "100100011",
       "001001000",
       "101101100",
       "001000000",
       "010000000",
       "001000000",
       "111110101",
       "011010001",
       "010001001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001001000",
       "011011010",
       "111111111",
       "100100011",
       "011010010",
       "111111111",
       "000000000",
       "110100100",
       "010000000",
       "111111110",
       "111110101",
       "010001000",
       "111110110",
       "111111111",
       "111111111",
       "111111111",
       "001001000",
       "001001000",
       "111111111",
       "100100011",
       "100011011",
       "111111110",
       "001000000",
       "111110101",
       "100011010",
       "111111110",
       "111110101",
       "101011011",
       "111110101",
       "111111111",
       "111111111",
       "111111111",
       "100010010",
       "100010010",
       "100011010",
       "100100011",
       "100100011",
       "110110101",
       "001000000",
       "111110110",
       "111111110",
       "111111110",
       "111110101",
       "101100100",
       "110101100",
       "111111111",
       "111111111",
       "111111111",
       "010001000",
       "011010001",
       "110101100",
       "100100011",
       "100100100",
       "110110101",
       "001000000",
       "001000000",
       "010001001",
       "111110110",
       "111111110",
       "011010001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011010",
       "010001000",
       "101100010",
       "100100011",
       "100100100",
       "101100100",
       "001001001",
       "001000000",
       "000000000",
       "100011011",
       "000000000",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "011001001",
       "101100011",
       "101100011",
       "100100011",
       "000000000",
       "100100011",
       "100011011",
       "001001000",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100011011",
       "000000000",
       "111110101",
       "110101100",
       "000000000",
       "011011010",
       "111111111",
       "100011011",
       "100011011",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "000000000",
       "111111110",
       "101101011",
       "001000000",
       "011011010",
       "111111110",
       "110101100",
       "111111110",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "000000000",
       "010010001",
       "110110100",
       "000000000",
       "000000000",
       "111111110",
       "111110101",
       "110101100",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "000000000",
       "010001000",
       "001000000",
       "001001001",
       "000000000",
       "011010001",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "001001001",
       "001001000",
       "001001010",
       "001001010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "000001000",
       "000001000",
       "000000001",
       "011011100",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "000000000",
       "111111111",
       "001001010",
       "010011100",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "001001001",
       "111111111",
       "000001001",
       "001010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010010",
       "010010010",
       "000000000",
       "111111111",
       "000001001",
       "001010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011011011",
       "011011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

