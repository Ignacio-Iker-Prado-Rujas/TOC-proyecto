------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : patron8b_100x100_color.ppm 
--- Filas    : 100 
--- Columnas : 100 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 8 bits
--- De cada palabra hay 3 bits para rojo y verde y 2 para azul: "RRRGGGBB" 256 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_8b_patron8b_100x100_color is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(14-1 downto 0);
    dout : out std_logic_vector(8-1 downto 0) 
  );
end ROM_RGB_8b_patron8b_100x100_color;


architecture BEHAVIORAL of ROM_RGB_8b_patron8b_100x100_color is
  signal addr_int  : natural range 0 to 2**14-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBB"
       "00111110",
       "11111111",
       "00111110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11111111",
       "11100100",
       "11111111",
       "00111110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11111111",
       "00111110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "00111101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11100100",
       "11100100",
       "11100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "01101101",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01101101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "10010011",
       "11111111",
       "10010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "00000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

