------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : game-over-negro.ppm 
--- Filas    : 34 
--- Columnas : 128 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_game-over-negro is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(13-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_game-over-negro;


architecture BEHAVIORAL of ROM_RGB_9b_game-over-negro is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100101",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101101100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "101101110",
       "101101101",
       "100100101",
       "111111111",
       "100100101",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "101101111",
       "101101110",
       "101101101",
       "111111111",
       "111111111",
       "101101110",
       "101101110",
       "101101110",
       "101101110",
       "111111111",
       "111111111",
       "101101110",
       "101101110",
       "100100110",
       "101101110",
       "111111111",
       "101101110",
       "101101110",
       "101101110",
       "101101110",
       "100100111",
       "011011110",
       "011011101",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100101",
       "111111111",
       "101101110",
       "101101110",
       "111111111",
       "100100100",
       "111111111",
       "101101110",
       "101101110",
       "101101111",
       "100100110",
       "111111111",
       "101101110",
       "101101110",
       "100101110",
       "101101110",
       "101101110",
       "101101110",
       "100100110",
       "101101110",
       "100101110",
       "100100101",
       "111111111",
       "101101101",
       "101101110",
       "101101110",
       "101101110",
       "100101110",
       "100100101",
       "111111111",
       "100100101",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "101101110",
       "111111111",
       "111111111",
       "100100110",
       "011011101",
       "011011101",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "101101111",
       "101101111",
       "100100101",
       "111111111",
       "100100101",
       "111111111",
       "100101110",
       "101101111",
       "101101110",
       "111111111",
       "111111111",
       "100101110",
       "100100110",
       "100100110",
       "111111111",
       "100100100",
       "111111111",
       "100101110",
       "101101110",
       "100100110",
       "011011110",
       "010010101",
       "010010100",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "101101110",
       "101101110",
       "100100110",
       "101101110",
       "111111111",
       "111111111",
       "101101110",
       "101101111",
       "101101111",
       "100100110",
       "111111111",
       "100100101",
       "100011110",
       "100100110",
       "111111111",
       "101101110",
       "100100110",
       "100011110",
       "100100110",
       "011011101",
       "011011101",
       "111111111",
       "111111111",
       "101101110",
       "101101110",
       "101101111",
       "111111111",
       "100100101",
       "011011100",
       "111111111",
       "100100101",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "101101110",
       "100100111",
       "111111111",
       "100100101",
       "111111111",
       "010011100",
       "010010101",
       "111111111",
       "000000000",
       "100100100",
       "111111111",
       "100100110",
       "100100110",
       "100100110",
       "111111111",
       "000000000",
       "111111111",
       "101101110",
       "101101111",
       "101101110",
       "111111111",
       "111111111",
       "100101110",
       "011100110",
       "011011110",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "100100110",
       "011011110",
       "111111111",
       "010010011",
       "010001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "101101111",
       "101101110",
       "111111111",
       "111111111",
       "100100110",
       "100100110",
       "111111111",
       "111111111",
       "100100110",
       "100100110",
       "011011110",
       "111111111",
       "111111111",
       "011011110",
       "111111111",
       "111111111",
       "100100110",
       "011100110",
       "011011110",
       "111111111",
       "011011101",
       "011010101",
       "111111111",
       "111111111",
       "100101110",
       "100100110",
       "100100110",
       "111111111",
       "011011110",
       "010010101",
       "010010100",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100110",
       "100100110",
       "111111111",
       "000000000",
       "111111111",
       "010010100",
       "010010101",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "100100110",
       "100100110",
       "011011110",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "101101111",
       "101101110",
       "111111111",
       "101101111",
       "011011101",
       "011011101",
       "010010101",
       "111111111",
       "000000000",
       "111111111",
       "011011101",
       "011100110",
       "010010101",
       "111111111",
       "111111111",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100101110",
       "100100110",
       "111111111",
       "111111111",
       "100100110",
       "100100110",
       "111111111",
       "111111111",
       "100100110",
       "011100101",
       "010011101",
       "111111111",
       "111111111",
       "011010101",
       "111111111",
       "111111111",
       "011100110",
       "011011101",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "111111111",
       "111111111",
       "100100110",
       "100100111",
       "011100110",
       "111111111",
       "010010101",
       "010010101",
       "010010100",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "100100110",
       "011011110",
       "111111111",
       "000000000",
       "100100100",
       "111111111",
       "010010101",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "100100101",
       "011011110",
       "011011110",
       "111111111",
       "100100100",
       "111111111",
       "100100101",
       "100100110",
       "100100110",
       "101101110",
       "011100110",
       "010011101",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "011011110",
       "010011101",
       "111111111",
       "111111111",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "100101111",
       "100100110",
       "111111111",
       "111111111",
       "100100110",
       "011100110",
       "111111111",
       "111111111",
       "011011110",
       "011011101",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "111111111",
       "111111111",
       "011011110",
       "010011101",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "111111111",
       "111111111",
       "011011101",
       "011011110",
       "011011110",
       "111111111",
       "010010101",
       "001010100",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "101101110",
       "100100110",
       "011011101",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "011100110",
       "111111111",
       "011011110",
       "011011110",
       "011011100",
       "111111111",
       "100100100",
       "111111111",
       "100100110",
       "100100110",
       "100100110",
       "011011110",
       "010010101",
       "010010100",
       "001010011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "001001010",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "101101110",
       "100100110",
       "100100110",
       "111111111",
       "111111111",
       "011011110",
       "011011110",
       "100100110",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "111111111",
       "111111111",
       "010011101",
       "010011101",
       "010010101",
       "111111111",
       "010010011",
       "111111111",
       "100100100",
       "111111111",
       "011100110",
       "011011110",
       "011011110",
       "111111111",
       "010010100",
       "001001011",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100101",
       "100100110",
       "011011101",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "011011101",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "111111111",
       "011011110",
       "011011110",
       "010011101",
       "111111111",
       "111111111",
       "100100110",
       "100100110",
       "100100111",
       "011100110",
       "011011110",
       "010010100",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011100110",
       "010010101",
       "111111111",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100110",
       "100100110",
       "011011110",
       "111111111",
       "111111111",
       "011011110",
       "011011110",
       "011011110",
       "111111111",
       "011011101",
       "010011101",
       "010010101",
       "111111111",
       "010011100",
       "111111111",
       "100100100",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "010010011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "011011110",
       "111111111",
       "010010011",
       "001001010",
       "001001001",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100110",
       "100100110",
       "011011110",
       "111111111",
       "000000000",
       "000000000",
       "100101100",
       "111111111",
       "100100100",
       "000000000",
       "111111111",
       "011011110",
       "111111111",
       "011011110",
       "011011110",
       "010011101",
       "111111111",
       "111111111",
       "100100110",
       "011100110",
       "011011110",
       "011011101",
       "010010101",
       "001001100",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "100100111",
       "011011110",
       "010011101",
       "111111111",
       "010001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100110",
       "100100111",
       "011011110",
       "111111111",
       "111111111",
       "011011110",
       "011011110",
       "011011101",
       "111111111",
       "011011101",
       "010011101",
       "010010101",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "011011110",
       "010011101",
       "111111111",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "011011110",
       "011011110",
       "111111111",
       "010010100",
       "001001010",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "100100110",
       "011100110",
       "011011110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "111111111",
       "011011110",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "011011101",
       "011011110",
       "011011110",
       "010011101",
       "010010100",
       "001001011",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "100011110",
       "011011110",
       "010011101",
       "010010011",
       "010001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011100110",
       "011100110",
       "011011110",
       "111111111",
       "111111111",
       "010011101",
       "010011110",
       "010010101",
       "111111111",
       "111111111",
       "010011101",
       "010010100",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010011101",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011100110",
       "010011101",
       "011011100",
       "010010100",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011100101",
       "011011110",
       "011011110",
       "111111111",
       "011011110",
       "011011110",
       "100100110",
       "100011101",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "011011101",
       "010011110",
       "010011110",
       "010010100",
       "001010100",
       "001001011",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "010010100",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011100110",
       "011011110",
       "011011101",
       "111111111",
       "111111111",
       "011011110",
       "010010101",
       "010010101",
       "111111111",
       "111111111",
       "010010101",
       "010010100",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "010010100",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "011011110",
       "011011110",
       "111111111",
       "010010100",
       "001010011",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "011011101",
       "111111111",
       "111111111",
       "011100101",
       "011011110",
       "011011110",
       "111111111",
       "100100100",
       "111111111",
       "011100101",
       "111111111",
       "011011110",
       "010011101",
       "010010101",
       "111111111",
       "111111111",
       "011010101",
       "010010101",
       "010010101",
       "010010100",
       "111111111",
       "001001100",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "010011110",
       "010011100",
       "111111111",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011011110",
       "011011111",
       "010011101",
       "111111111",
       "111111111",
       "010010101",
       "010010101",
       "010010101",
       "111111111",
       "111111111",
       "010010101",
       "010010100",
       "010010100",
       "010010011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "100100110",
       "011100110",
       "011011101",
       "111111111",
       "010010100",
       "001010100",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011011101",
       "010011110",
       "011011101",
       "111111111",
       "111111111",
       "011011110",
       "011011111",
       "011011101",
       "111111111",
       "111111111",
       "100011101",
       "111111111",
       "111111111",
       "011100110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "011010101",
       "111111111",
       "010011101",
       "010010100",
       "111111111",
       "010001100",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "010011110",
       "010010100",
       "111111111",
       "010010011",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "011011101",
       "010011110",
       "011011101",
       "111111111",
       "111111111",
       "010010100",
       "010010100",
       "010010100",
       "111111111",
       "111111111",
       "010010100",
       "001010100",
       "001001011",
       "001010010",
       "111111111",
       "000000000",
       "111111111",
       "011011101",
       "011011110",
       "010010101",
       "111111111",
       "010010100",
       "111111111",
       "100100100",
       "111111111",
       "100100110",
       "011011110",
       "011011110",
       "111111111",
       "010010101",
       "001010100",
       "010010011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010011100",
       "010011110",
       "010010101",
       "111111111",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "011011110",
       "111111111",
       "100100101",
       "011011101",
       "011011111",
       "011011110",
       "111111111",
       "111111111",
       "011011101",
       "111111111",
       "010011110",
       "010010101",
       "111111111",
       "010010100",
       "010010011",
       "001010011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "001001011",
       "010010010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010011100",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "001010100",
       "010010011",
       "111111111",
       "111111111",
       "010010100",
       "001010100",
       "001010100",
       "111111111",
       "100100100",
       "000000000",
       "111111111",
       "011100110",
       "011011110",
       "010010101",
       "111111111",
       "010010011",
       "011011101",
       "111111111",
       "111111111",
       "100100110",
       "011100111",
       "011011110",
       "111111111",
       "010010100",
       "010010100",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "010010101",
       "010010100",
       "111111111",
       "111111111",
       "010010101",
       "010010101",
       "010010101",
       "111111111",
       "111111111",
       "011010101",
       "111111111",
       "111111111",
       "011100101",
       "011011111",
       "010011110",
       "011011101",
       "111111111",
       "011011101",
       "111111111",
       "010010101",
       "010010101",
       "111111111",
       "010010100",
       "001010011",
       "010010100",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "010011110",
       "010010101",
       "111111111",
       "111111111",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "010011101",
       "010010101",
       "111111111",
       "111111111",
       "010010100",
       "001001011",
       "111111111",
       "100100100",
       "111111111",
       "001001011",
       "001010011",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010101",
       "111111111",
       "111111111",
       "010010101",
       "111111111",
       "111111111",
       "011100110",
       "011011110",
       "011011110",
       "111111111",
       "010010100",
       "010010100",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010010100",
       "010010100",
       "111111111",
       "111111111",
       "010010100",
       "001001011",
       "001001100",
       "111111111",
       "111111111",
       "010010101",
       "111111111",
       "100100100",
       "111111111",
       "010010101",
       "010010101",
       "011011101",
       "111111111",
       "010010101",
       "111111111",
       "010011101",
       "001010011",
       "111111111",
       "010010100",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "011011110",
       "010011101",
       "010010100",
       "111111111",
       "111111111",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010010101",
       "010010100",
       "111111111",
       "111111111",
       "001001011",
       "001001010",
       "111111111",
       "000000000",
       "111111111",
       "001001011",
       "001010011",
       "001001011",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "011011110",
       "011011110",
       "010010100",
       "111111111",
       "111111111",
       "010010101",
       "111111111",
       "111111111",
       "011011101",
       "010010101",
       "010010101",
       "111111111",
       "010010100",
       "001001010",
       "001001010",
       "111111111",
       "101101101",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010010100",
       "010010011",
       "111111111",
       "111111111",
       "010010100",
       "001001010",
       "001001011",
       "111111111",
       "111111111",
       "010010101",
       "111111111",
       "100100100",
       "111111111",
       "010011101",
       "010010100",
       "010010100",
       "111111111",
       "010001100",
       "111111111",
       "001001011",
       "010010011",
       "111111111",
       "001001011",
       "001001010",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "010010101",
       "010011101",
       "010010100",
       "111111111",
       "010010011",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "010010100",
       "010010100",
       "111111111",
       "111111111",
       "001001010",
       "001001010",
       "111111111",
       "000000000",
       "100100101",
       "111111111",
       "001001011",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "111111111",
       "011011101",
       "010010101",
       "010010100",
       "111111111",
       "010010011",
       "010010100",
       "111111111",
       "111111111",
       "010010100",
       "010010100",
       "001010100",
       "111111111",
       "001001010",
       "001001010",
       "000001010",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "010010011",
       "111111111",
       "111111111",
       "001001010",
       "001001010",
       "111111111",
       "111111111",
       "010010011",
       "010010100",
       "111111111",
       "111111111",
       "010010100",
       "001001011",
       "001010100",
       "010010011",
       "001001010",
       "001001011",
       "001001010",
       "001001011",
       "111111111",
       "111111111",
       "001001010",
       "001001010",
       "001001011",
       "111111111",
       "100100100",
       "111111111",
       "010010100",
       "001001011",
       "001001011",
       "111111111",
       "001001011",
       "001001010",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100101",
       "111111111",
       "001010011",
       "001010010",
       "001001010",
       "001001001",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "111111111",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "100100100",
       "111111111",
       "010010100",
       "010010100",
       "001001011",
       "111111111",
       "001001011",
       "001001011",
       "111111111",
       "111111111",
       "010010011",
       "001001011",
       "001001011",
       "111111111",
       "001001010",
       "000001001",
       "000000001",
       "001000001",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100101",
       "111111111",
       "001001010",
       "001001010",
       "111111111",
       "111111111",
       "100100101",
       "111111111",
       "001001010",
       "001001011",
       "001001011",
       "111111111",
       "001001011",
       "001001010",
       "000000010",
       "000000001",
       "000000001",
       "000000001",
       "000000001",
       "000000001",
       "111111111",
       "111111111",
       "000000010",
       "000001010",
       "000001010",
       "001001001",
       "111111111",
       "001001010",
       "001001011",
       "000001011",
       "000001001",
       "000001001",
       "001000011",
       "000001001",
       "111111111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100101",
       "111111111",
       "001001010",
       "001001010",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "111111111",
       "001001011",
       "001001011",
       "111111111",
       "000000000",
       "111111111",
       "010010011",
       "010010100",
       "001001011",
       "000001010",
       "001001001",
       "001001011",
       "000001001",
       "111111111",
       "001001010",
       "001001010",
       "000001011",
       "000001001",
       "001000001",
       "111111111",
       "000000001",
       "000000001",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "101101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101101101",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "100100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101101101",
       "111111111",
       "111111111",
       "100100100",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

