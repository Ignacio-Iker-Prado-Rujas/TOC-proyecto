--------------------------------------------------------------------------------
-- Felipe Machado Sanchez
-- Departameto de Tecnologia Electronica
-- Universidad Rey Juan Carlos
-- http://gtebim.es/~fmachado
--
-- ROM para los caractere ASCII, solo estan los caracteres alfanumericos
-- y alguno mas, como lo dos puntos, comas,...
-- las minusculas estan en mayusculas, asi que hay dos A, dos B,...


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;

entity romchar is
  generic (
    gbitsprofBRAM       : natural := 11; -- 2048 posiciones
    gbitsBRAM           : natural := 8  -- palabra de 8 bits
  );
  port(
    clka         : in std_logic;
    addra        : in std_logic_vector(gbitsprofBRAM-1 downto 0);
    douta        : out std_logic_vector(gbitsBRAM-1 downto 0)
  );
end romchar;

architecture BEHAVIOURAL of romchar is

  signal addra_int   : natural range 0 to 2**gbitsprofBRAM-1;

  type  memostruct is array (natural range<>) of std_logic_vector(gbitsBRAM-1 downto 0);
 
  constant datosChar : memostruct := (
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "01101110", "01110110",
            "01100110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00011000", "00011000", "00111000", "00011000",
            "00011000", "00011000", "01111110", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "00000110", "00001100",
            "00110000", "01100000", "01111110", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "00000110", "00011100",
            "00000110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000110", "00001110", "00011110", "01100110",
            "01111111", "00000110", "00000110", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "01111110", "01100000", "01111100", "00000110",
            "00000110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "01100000", "01111100",
            "01100110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "01111110", "01100110", "00001100", "00011000",
            "00011000", "00011000", "00011000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "01100110", "00111100",
            "01100110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00111100", "01100110", "01100110", "00111110",
            "00000110", "01100110", "00111100", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00011000", "00011000", "00000000",
            "00011000", "00011000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00011000", "00011000", "00000000",
            "00011000", "00011000", "00001000", "00010000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00001100", "00011000", "00110000",
            "01100000", "00110000", "00011000", "00001100",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "11111111",
            "00000000", "11111111", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00110000", "00011000", "00001100",
            "00000110", "00001100", "00011000", "00110000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01000110",
            "00000110", "00000110", "00001100", "00011000",
            "00110000", "00000000", "00110000", "00110000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01101110", "01101110", "01100000", "01100010",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011000", "00111100",
            "01100110", "01111110", "01100110", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111100", "01100110",
            "01100110", "01111100", "01100110", "01100110",
            "01111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100000", "01100000", "01100000", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111000", "01101100",
            "01100110", "01100110", "01100110", "01101100",
            "01111000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "01100000",
            "01100000", "01111000", "01100000", "01100000",
            "01111110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "01100000",
            "01100000", "01111000", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100000", "01101110", "01100110", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "01100110", "01111110", "01100110", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "00011000",
            "00011000", "00011000", "00011000", "00011000",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011110", "00001100",
            "00001100", "00001100", "00001100", "01101100",
            "00111000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01101100",
            "01111000", "01110000", "01111000", "01101100",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100000", "01100000",
            "01100000", "01100000", "01100000", "01100000",
            "01111110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100011", "01110111",
            "01111111", "01101011", "01100011", "01100011",
            "01100011", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01110110",
            "01111110", "01111110", "01101110", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100110", "01100110", "01100110", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111100", "01100110",
            "01100110", "01111100", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100110", "01100110", "01100110", "00111100",
            "00001110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111100", "01100110",
            "01100110", "01111100", "01111000", "01101100",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100000", "00111100", "00000110", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "00011000",
            "00011000", "00011000", "00011000", "00011000",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "01100110", "01100110", "01100110", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "01100110", "01100110", "01100110", "00111100",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100011", "01100011",
            "01100011", "01101011", "01111111", "01110111",
            "01100011", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "00111100", "00011000", "00111100", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "01100110", "00111100", "00011000", "00011000",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "00000110",
            "00001100", "00011000", "00110000", "01100000",
            "01111110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "00110000",
            "00110000", "00110000", "00110000", "00110000",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011000", "00011000",
            "00011000", "00011000", "01111110", "00111100",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "00001100",
            "00001100", "00001100", "00001100", "00001100",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00011000",
            "00111100", "01111110", "00011000", "00011000",
            "00011000", "00011000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00010000",
            "00110000", "01111111", "01111111", "00110000",
            "00010000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011000", "00011000",
            "00011000", "00011000", "00000000", "00000000",
            "00011000", "00000000", "01100110", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100110", "01100110",
            "11111111", "01100110", "11111111", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011000", "00111110",
            "01100000", "00111100", "00000110", "01111100",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100010", "01100110",
            "00001100", "00011000", "00110000", "01100110",
            "01000110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "00111100", "00111000", "01100111", "01100110",
            "00111111", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000110", "00001100",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00001100", "00011000",
            "00110000", "00110000", "00110000", "00011000",
            "00001100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00110000", "00011000",
            "00001100", "00001100", "00001100", "00011000",
            "00110000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "01100110",
            "00111100", "11111111", "00111100", "01100110",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00011000",
            "00011000", "01111110", "00011000", "00011000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00011000",
            "00011000", "00110000", "00000000", "00000000",
            "00000000", "01111110", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00011000",
            "00011000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000011",
            "00000110", "00001100", "00011000", "00110000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00011000", "00111100",
            "01100110", "01111110", "01100110", "01100110",
            "01100110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111100", "01100110",
            "01100110", "01111100", "01100110", "01100110",
            "01111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00111100", "01100110",
            "01100000", "01100000", "01100000", "01100110",
            "00111100", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111000", "01101100",
            "01100110", "01100110", "01100110", "01101100",
            "01111000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "01100000",
            "01100000", "01111000", "01100000", "01100000",
            "01111110", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111110", "01100000",
            "01100000", "01111000", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01111000", "01100000",
            "01100000", "01100000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "01111000",
            "01111000", "01111000", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "01100000", "01100000",
            "01100000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000",
            "00000000", "00000000", "00000000", "00000000"
            );

begin 

 addra_int <= TO_INTEGER(unsigned(addra));

  P: process (clka)
  begin
    if clka'event and clka='1' then
      douta <= datosChar(addra_int);
    end if;
  end process;

end BEHAVIOURAL;
